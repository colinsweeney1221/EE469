module lab1 (out, in);
	output out;
	input in;
	
	assign out = in;
	
endmodule