module control();
endmodule
