module lab2 (out, in);
	output out;
	input in;
	
	assign out = in;
	
endmodule